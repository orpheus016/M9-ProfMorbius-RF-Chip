magic
tech gf180mcuD
magscale 1 10
timestamp 1758388245
<< nwell >>
rect -2080 -120 -536 452
rect -60 -120 1484 452
rect -7740 -1480 -6162 -964
rect 5380 -1480 6958 -964
rect 5940 -2740 6494 -2304
<< pwell >>
rect -5440 -1020 -3064 -640
rect -2980 -1020 -604 -640
rect -20 -1020 2356 -640
rect 2480 -1020 4856 -640
rect -5440 -1460 -824 -1080
rect 240 -1380 4856 -1080
rect 204 -1460 4856 -1380
rect -6780 -2200 -3284 -1920
rect -7440 -5440 -6768 -3224
rect -6580 -31940 -5908 -3224
rect -5780 -31940 -5108 -3224
rect -4980 -31940 -4308 -3224
rect -4180 -31940 -3508 -3224
rect -2580 -31940 -1908 -3224
rect -1780 -31940 -1108 -3224
rect 420 -31940 1092 -3224
rect 1220 -31940 1892 -3224
rect 2020 -31940 2692 -3224
rect 2820 -31940 3492 -3224
rect 3620 -31940 4292 -3224
rect 5220 -31940 5892 -3224
rect 6040 -3340 6430 -3028
rect -2380 -32080 -2100 -32076
rect -1580 -32080 -1300 -32076
rect -6480 -33000 -6100 -32080
rect -5680 -33000 -5300 -32080
rect -4880 -33000 -4500 -32080
rect -4080 -32100 -3780 -32080
rect -2280 -32100 -2100 -32080
rect -4080 -33000 -3700 -32100
rect -2480 -33820 -2100 -32100
rect -1680 -33820 -1300 -32080
rect 620 -32140 900 -32084
rect 1420 -32140 1700 -32084
rect 2220 -32140 2500 -32084
rect 3020 -32140 3300 -32084
rect 620 -32780 1000 -32140
rect 1420 -32780 1800 -32140
rect 2220 -32780 2600 -32140
rect 3020 -32780 3400 -32140
rect 3820 -32780 4200 -32084
rect 5420 -32380 5800 -32076
rect -6580 -62640 -5908 -33924
rect -5780 -62640 -5108 -33924
rect -4980 -62640 -4308 -33924
rect -4180 -62640 -3508 -33924
rect -2580 -62640 -1908 -33924
rect -1780 -62640 -1108 -33924
rect 420 -62600 1092 -33884
rect 1220 -62600 1892 -33884
rect 2020 -62600 2692 -33884
rect 2820 -62600 3492 -33884
rect 3620 -62600 4292 -33884
rect 5220 -62600 5892 -33884
<< nmos >>
rect -5372 -808 -3132 -752
rect -2912 -808 -672 -752
rect 48 -808 2288 -752
rect 2548 -808 4788 -752
rect -5372 -1248 -892 -1192
rect 308 -1248 4788 -1192
rect -6712 -2088 -3352 -2032
rect -6712 -2468 -3352 -2412
rect 6262 -3272 6318 -3096
rect -6268 -32932 -6212 -32148
rect -5468 -32932 -5412 -32148
rect -4668 -32932 -4612 -32148
rect -3868 -32932 -3812 -32148
rect -2268 -33712 -2212 -32144
rect -1468 -33712 -1412 -32144
rect 732 -32712 788 -32152
rect 1532 -32712 1588 -32152
rect 2332 -32712 2388 -32152
rect 3132 -32712 3188 -32152
rect 3932 -32712 3988 -32152
rect 5532 -32312 5588 -32144
<< pmos >>
rect 6264 -2610 6320 -2434
<< ndiff >>
rect -5372 -677 -3132 -664
rect -5372 -723 -5359 -677
rect -3145 -723 -3132 -677
rect -5372 -752 -3132 -723
rect -2912 -677 -672 -664
rect -2912 -723 -2899 -677
rect -685 -723 -672 -677
rect 48 -677 2288 -664
rect -2912 -752 -672 -723
rect -5372 -837 -3132 -808
rect -5372 -883 -5359 -837
rect -3145 -883 -3132 -837
rect -5372 -896 -3132 -883
rect -2912 -837 -672 -808
rect -2912 -883 -2899 -837
rect -685 -883 -672 -837
rect 48 -723 61 -677
rect 2275 -723 2288 -677
rect 48 -752 2288 -723
rect 2548 -677 4788 -664
rect 2548 -723 2561 -677
rect 4775 -723 4788 -677
rect 2548 -752 4788 -723
rect 48 -837 2288 -808
rect -2912 -896 -672 -883
rect 48 -883 61 -837
rect 2275 -883 2288 -837
rect 48 -896 2288 -883
rect 2548 -837 4788 -808
rect 2548 -883 2561 -837
rect 4775 -883 4788 -837
rect 2548 -896 4788 -883
rect -5372 -1117 -892 -1104
rect -5372 -1163 -5359 -1117
rect -905 -1163 -892 -1117
rect -5372 -1192 -892 -1163
rect 308 -1117 4788 -1104
rect 308 -1163 321 -1117
rect 4775 -1163 4788 -1117
rect 308 -1192 4788 -1163
rect -5372 -1277 -892 -1248
rect -5372 -1323 -5359 -1277
rect -905 -1323 -892 -1277
rect -5372 -1336 -892 -1323
rect 308 -1277 4788 -1248
rect 308 -1323 321 -1277
rect 4775 -1323 4788 -1277
rect 308 -1336 4788 -1323
rect -6712 -1957 -3352 -1944
rect -6712 -2003 -6699 -1957
rect -3365 -2003 -3352 -1957
rect -6712 -2032 -3352 -2003
rect -6712 -2117 -3352 -2088
rect -6712 -2163 -6699 -2117
rect -3365 -2163 -3352 -2117
rect -6712 -2176 -3352 -2163
rect -6712 -2337 -3352 -2324
rect -6712 -2383 -6699 -2337
rect -3365 -2383 -3352 -2337
rect -6712 -2412 -3352 -2383
rect -6712 -2497 -3352 -2468
rect -6712 -2543 -6699 -2497
rect -3365 -2543 -3352 -2497
rect -6712 -2556 -3352 -2543
rect 6174 -3109 6262 -3096
rect 6174 -3259 6187 -3109
rect 6233 -3259 6262 -3109
rect 6174 -3272 6262 -3259
rect 6318 -3109 6406 -3096
rect 6318 -3259 6347 -3109
rect 6393 -3259 6406 -3109
rect 6318 -3272 6406 -3259
rect -6356 -32161 -6268 -32148
rect -6356 -32919 -6343 -32161
rect -6297 -32919 -6268 -32161
rect -6356 -32932 -6268 -32919
rect -6212 -32161 -6124 -32148
rect -6212 -32919 -6183 -32161
rect -6137 -32919 -6124 -32161
rect -6212 -32932 -6124 -32919
rect -5556 -32161 -5468 -32148
rect -5556 -32919 -5543 -32161
rect -5497 -32919 -5468 -32161
rect -5556 -32932 -5468 -32919
rect -5412 -32161 -5324 -32148
rect -5412 -32919 -5383 -32161
rect -5337 -32919 -5324 -32161
rect -5412 -32932 -5324 -32919
rect -4756 -32161 -4668 -32148
rect -4756 -32919 -4743 -32161
rect -4697 -32919 -4668 -32161
rect -4756 -32932 -4668 -32919
rect -4612 -32161 -4524 -32148
rect -4612 -32919 -4583 -32161
rect -4537 -32919 -4524 -32161
rect -4612 -32932 -4524 -32919
rect -3956 -32161 -3868 -32148
rect -3956 -32919 -3943 -32161
rect -3897 -32919 -3868 -32161
rect -3956 -32932 -3868 -32919
rect -3812 -32161 -3724 -32148
rect -3812 -32919 -3783 -32161
rect -3737 -32919 -3724 -32161
rect -3812 -32932 -3724 -32919
rect -2356 -32157 -2268 -32144
rect -2356 -33699 -2343 -32157
rect -2297 -33699 -2268 -32157
rect -2356 -33712 -2268 -33699
rect -2212 -32157 -2124 -32144
rect -2212 -33699 -2183 -32157
rect -2137 -33699 -2124 -32157
rect -2212 -33712 -2124 -33699
rect -1556 -32157 -1468 -32144
rect -1556 -33699 -1543 -32157
rect -1497 -33699 -1468 -32157
rect -1556 -33712 -1468 -33699
rect -1412 -32157 -1324 -32144
rect -1412 -33699 -1383 -32157
rect -1337 -33699 -1324 -32157
rect 644 -32165 732 -32152
rect 644 -32699 657 -32165
rect 703 -32699 732 -32165
rect 644 -32712 732 -32699
rect 788 -32165 876 -32152
rect 788 -32699 817 -32165
rect 863 -32699 876 -32165
rect 788 -32712 876 -32699
rect 1444 -32165 1532 -32152
rect 1444 -32699 1457 -32165
rect 1503 -32699 1532 -32165
rect 1444 -32712 1532 -32699
rect 1588 -32165 1676 -32152
rect 1588 -32699 1617 -32165
rect 1663 -32699 1676 -32165
rect 1588 -32712 1676 -32699
rect 2244 -32165 2332 -32152
rect 2244 -32699 2257 -32165
rect 2303 -32699 2332 -32165
rect 2244 -32712 2332 -32699
rect 2388 -32165 2476 -32152
rect 2388 -32699 2417 -32165
rect 2463 -32699 2476 -32165
rect 2388 -32712 2476 -32699
rect 3044 -32165 3132 -32152
rect 3044 -32699 3057 -32165
rect 3103 -32699 3132 -32165
rect 3044 -32712 3132 -32699
rect 3188 -32165 3276 -32152
rect 3188 -32699 3217 -32165
rect 3263 -32699 3276 -32165
rect 3188 -32712 3276 -32699
rect 3844 -32165 3932 -32152
rect 3844 -32699 3857 -32165
rect 3903 -32699 3932 -32165
rect 3844 -32712 3932 -32699
rect 3988 -32165 4076 -32152
rect 3988 -32699 4017 -32165
rect 4063 -32699 4076 -32165
rect 5444 -32157 5532 -32144
rect 5444 -32299 5457 -32157
rect 5503 -32299 5532 -32157
rect 5444 -32312 5532 -32299
rect 5588 -32157 5676 -32144
rect 5588 -32299 5617 -32157
rect 5663 -32299 5676 -32157
rect 5588 -32312 5676 -32299
rect 3988 -32712 4076 -32699
rect -1412 -33712 -1324 -33699
<< pdiff >>
rect -1894 253 -1768 266
rect -1894 79 -1881 253
rect -1835 79 -1768 253
rect -1894 66 -1768 79
rect -848 253 -722 266
rect -848 79 -781 253
rect -735 79 -722 253
rect -848 66 -722 79
rect 126 253 252 266
rect 126 79 139 253
rect 185 79 252 253
rect 126 66 252 79
rect 1172 253 1298 266
rect 1172 79 1239 253
rect 1285 79 1298 253
rect 1172 66 1298 79
rect 6176 -2447 6264 -2434
rect 6176 -2597 6189 -2447
rect 6235 -2597 6264 -2447
rect 6176 -2610 6264 -2597
rect 6320 -2447 6408 -2434
rect 6320 -2597 6349 -2447
rect 6395 -2597 6408 -2447
rect 6320 -2610 6408 -2597
<< ndiffc >>
rect -5359 -723 -3145 -677
rect -2899 -723 -685 -677
rect -5359 -883 -3145 -837
rect -2899 -883 -685 -837
rect 61 -723 2275 -677
rect 2561 -723 4775 -677
rect 61 -883 2275 -837
rect 2561 -883 4775 -837
rect -5359 -1163 -905 -1117
rect 321 -1163 4775 -1117
rect -5359 -1323 -905 -1277
rect 321 -1323 4775 -1277
rect -6699 -2003 -3365 -1957
rect -6699 -2163 -3365 -2117
rect -6699 -2383 -3365 -2337
rect -6699 -2543 -3365 -2497
rect 6187 -3259 6233 -3109
rect 6347 -3259 6393 -3109
rect -6343 -32919 -6297 -32161
rect -6183 -32919 -6137 -32161
rect -5543 -32919 -5497 -32161
rect -5383 -32919 -5337 -32161
rect -4743 -32919 -4697 -32161
rect -4583 -32919 -4537 -32161
rect -3943 -32919 -3897 -32161
rect -3783 -32919 -3737 -32161
rect -2343 -33699 -2297 -32157
rect -2183 -33699 -2137 -32157
rect -1543 -33699 -1497 -32157
rect -1383 -33699 -1337 -32157
rect 657 -32699 703 -32165
rect 817 -32699 863 -32165
rect 1457 -32699 1503 -32165
rect 1617 -32699 1663 -32165
rect 2257 -32699 2303 -32165
rect 2417 -32699 2463 -32165
rect 3057 -32699 3103 -32165
rect 3217 -32699 3263 -32165
rect 3857 -32699 3903 -32165
rect 4017 -32699 4063 -32165
rect 5457 -32299 5503 -32157
rect 5617 -32299 5663 -32157
<< pdiffc >>
rect -1881 79 -1835 253
rect -781 79 -735 253
rect 139 79 185 253
rect 1239 79 1285 253
rect 6189 -2597 6235 -2447
rect 6349 -2597 6395 -2447
<< psubdiff >>
rect -5372 -934 -3132 -896
rect -5372 -980 -5300 -934
rect -3160 -980 -3132 -934
rect -5372 -1000 -3132 -980
rect -2912 -934 -672 -896
rect -2912 -980 -2884 -934
rect -744 -980 -672 -934
rect -2912 -1000 -672 -980
rect 48 -934 2288 -896
rect 48 -980 120 -934
rect 2260 -980 2288 -934
rect 48 -1000 2288 -980
rect 2548 -934 4788 -896
rect 2548 -980 2576 -934
rect 4716 -980 4788 -934
rect 2548 -1000 4788 -980
rect -5372 -1374 -892 -1336
rect -5372 -1420 -5300 -1374
rect -905 -1420 -892 -1374
rect -5372 -1440 -892 -1420
rect 308 -1374 4788 -1336
rect 308 -1420 321 -1374
rect 4716 -1420 4788 -1374
rect 308 -1440 4788 -1420
rect -6712 -2227 -3352 -2176
rect -6712 -2273 -6660 -2227
rect -3380 -2273 -3352 -2227
rect -6712 -2324 -3352 -2273
rect 6064 -3109 6174 -3096
rect -7416 -3320 -6792 -3248
rect -7416 -5344 -7344 -3320
rect -6864 -5344 -6792 -3320
rect -7416 -5416 -6792 -5344
rect -6556 -3320 -5932 -3248
rect -6556 -31844 -6484 -3320
rect -6004 -31844 -5932 -3320
rect -6556 -31916 -5932 -31844
rect -5756 -3320 -5132 -3248
rect -5756 -31844 -5684 -3320
rect -5204 -31844 -5132 -3320
rect -5756 -31916 -5132 -31844
rect -4956 -3320 -4332 -3248
rect -4956 -31844 -4884 -3320
rect -4404 -31844 -4332 -3320
rect -4956 -31916 -4332 -31844
rect -4156 -3320 -3532 -3248
rect -4156 -31844 -4084 -3320
rect -3604 -31844 -3532 -3320
rect -4156 -31916 -3532 -31844
rect -2556 -3320 -1932 -3248
rect -2556 -31844 -2484 -3320
rect -2004 -31844 -1932 -3320
rect -2556 -31916 -1932 -31844
rect -1756 -3320 -1132 -3248
rect -1756 -31844 -1684 -3320
rect -1204 -31844 -1132 -3320
rect -1756 -31916 -1132 -31844
rect 444 -3320 1068 -3248
rect 444 -31844 516 -3320
rect 996 -31844 1068 -3320
rect 444 -31916 1068 -31844
rect 1244 -3320 1868 -3248
rect 1244 -31844 1316 -3320
rect 1796 -31844 1868 -3320
rect 1244 -31916 1868 -31844
rect 2044 -3320 2668 -3248
rect 2044 -31844 2116 -3320
rect 2596 -31844 2668 -3320
rect 2044 -31916 2668 -31844
rect 2844 -3320 3468 -3248
rect 2844 -31844 2916 -3320
rect 3396 -31844 3468 -3320
rect 2844 -31916 3468 -31844
rect 3644 -3320 4268 -3248
rect 3644 -31844 3716 -3320
rect 4196 -31844 4268 -3320
rect 3644 -31916 4268 -31844
rect 5244 -3320 5868 -3248
rect 6064 -3259 6084 -3109
rect 6130 -3259 6174 -3109
rect 6064 -3272 6174 -3259
rect 5244 -31844 5316 -3320
rect 5796 -31844 5868 -3320
rect 5244 -31916 5868 -31844
rect -6460 -32220 -6356 -32148
rect -6460 -32919 -6440 -32220
rect -6394 -32919 -6356 -32220
rect -6460 -32932 -6356 -32919
rect -5660 -32220 -5556 -32148
rect -5660 -32919 -5640 -32220
rect -5594 -32919 -5556 -32220
rect -5660 -32932 -5556 -32919
rect -4860 -32220 -4756 -32148
rect -4860 -32919 -4840 -32220
rect -4794 -32919 -4756 -32220
rect -4860 -32932 -4756 -32919
rect -4060 -32220 -3956 -32148
rect -4060 -32919 -4040 -32220
rect -3994 -32919 -3956 -32220
rect -4060 -32932 -3956 -32919
rect -2460 -32220 -2356 -32144
rect -2460 -33699 -2446 -32220
rect -2400 -33699 -2356 -32220
rect -2460 -33712 -2356 -33699
rect -1660 -32220 -1556 -32144
rect -1660 -33699 -1646 -32220
rect -1600 -33699 -1556 -32220
rect -1660 -33712 -1556 -33699
rect 876 -32220 980 -32152
rect 876 -32699 920 -32220
rect 966 -32699 980 -32220
rect 876 -32712 980 -32699
rect 1676 -32220 1780 -32152
rect 1676 -32699 1720 -32220
rect 1766 -32699 1780 -32220
rect 1676 -32712 1780 -32699
rect 2476 -32220 2580 -32152
rect 2476 -32699 2520 -32220
rect 2566 -32699 2580 -32220
rect 2476 -32712 2580 -32699
rect 3276 -32220 3380 -32152
rect 3276 -32699 3320 -32220
rect 3366 -32699 3380 -32220
rect 3276 -32712 3380 -32699
rect 4076 -32220 4180 -32152
rect 4076 -32699 4120 -32220
rect 4166 -32699 4180 -32220
rect 5676 -32211 5780 -32144
rect 5676 -32299 5720 -32211
rect 5766 -32299 5780 -32211
rect 5676 -32312 5780 -32299
rect 4076 -32712 4180 -32699
rect -6556 -34020 -5932 -33948
rect -6556 -62544 -6484 -34020
rect -6004 -62544 -5932 -34020
rect -6556 -62616 -5932 -62544
rect -5756 -34020 -5132 -33948
rect -5756 -62544 -5684 -34020
rect -5204 -62544 -5132 -34020
rect -5756 -62616 -5132 -62544
rect -4956 -34020 -4332 -33948
rect -4956 -62544 -4884 -34020
rect -4404 -62544 -4332 -34020
rect -4956 -62616 -4332 -62544
rect -4156 -34020 -3532 -33948
rect -4156 -62544 -4084 -34020
rect -3604 -62544 -3532 -34020
rect -4156 -62616 -3532 -62544
rect -2556 -34020 -1932 -33948
rect -2556 -62544 -2484 -34020
rect -2004 -62544 -1932 -34020
rect -2556 -62616 -1932 -62544
rect -1756 -34020 -1132 -33948
rect -1756 -62544 -1684 -34020
rect -1204 -62544 -1132 -34020
rect -1756 -62616 -1132 -62544
rect 444 -33980 1068 -33908
rect 444 -62504 516 -33980
rect 996 -62504 1068 -33980
rect 444 -62576 1068 -62504
rect 1244 -33980 1868 -33908
rect 1244 -62504 1316 -33980
rect 1796 -62504 1868 -33980
rect 1244 -62576 1868 -62504
rect 2044 -33980 2668 -33908
rect 2044 -62504 2116 -33980
rect 2596 -62504 2668 -33980
rect 2044 -62576 2668 -62504
rect 2844 -33980 3468 -33908
rect 2844 -62504 2916 -33980
rect 3396 -62504 3468 -33980
rect 2844 -62576 3468 -62504
rect 3644 -33980 4268 -33908
rect 3644 -62504 3716 -33980
rect 4196 -62504 4268 -33980
rect 3644 -62576 4268 -62504
rect 5244 -33980 5868 -33908
rect 5244 -62504 5316 -33980
rect 5796 -62504 5868 -33980
rect 5244 -62576 5868 -62504
<< nsubdiff >>
rect -2056 356 -560 428
rect -2056 -24 -1984 356
rect -632 -24 -560 356
rect -2056 -96 -560 -24
rect -36 356 1460 428
rect -36 -24 36 356
rect 1388 -24 1460 356
rect -36 -96 1460 -24
rect -7716 -1060 -6186 -988
rect -7716 -1384 -7644 -1060
rect -6258 -1384 -6186 -1060
rect 5404 -1060 6934 -988
rect -7716 -1456 -6186 -1384
rect 5404 -1384 5476 -1060
rect 6862 -1384 6934 -1060
rect 5404 -1456 6934 -1384
rect 6066 -2447 6176 -2434
rect 6066 -2597 6085 -2447
rect 6131 -2597 6176 -2447
rect 6066 -2610 6176 -2597
<< psubdiffcont >>
rect -5300 -980 -3160 -934
rect -2884 -980 -744 -934
rect 120 -980 2260 -934
rect 2576 -980 4716 -934
rect -5300 -1420 -905 -1374
rect 321 -1420 4716 -1374
rect -6660 -2273 -3380 -2227
rect 6084 -3259 6130 -3109
rect -6440 -32919 -6394 -32220
rect -5640 -32919 -5594 -32220
rect -4840 -32919 -4794 -32220
rect -4040 -32919 -3994 -32220
rect -2446 -33699 -2400 -32220
rect -1646 -33699 -1600 -32220
rect 920 -32699 966 -32220
rect 1720 -32699 1766 -32220
rect 2520 -32699 2566 -32220
rect 3320 -32699 3366 -32220
rect 4120 -32699 4166 -32220
rect 5720 -32299 5766 -32211
<< nsubdiffcont >>
rect 6085 -2597 6131 -2447
<< polysilicon >>
rect -5600 -740 -5480 -720
rect -5600 -820 -5580 -740
rect -5500 -760 -5480 -740
rect -540 -740 -420 -720
rect -5416 -760 -5372 -752
rect -5500 -800 -5372 -760
rect -5500 -820 -5480 -800
rect -5416 -808 -5372 -800
rect -3132 -808 -3088 -752
rect -2956 -808 -2912 -752
rect -672 -760 -628 -752
rect -540 -760 -520 -740
rect -672 -800 -520 -760
rect -672 -808 -628 -800
rect -5600 -840 -5480 -820
rect -540 -820 -520 -800
rect -440 -820 -420 -740
rect -540 -840 -420 -820
rect -180 -740 -60 -720
rect -180 -820 -160 -740
rect -80 -760 -60 -740
rect 4900 -740 5020 -720
rect 4 -760 48 -752
rect -80 -800 48 -760
rect -80 -820 -60 -800
rect 4 -808 48 -800
rect 2288 -808 2332 -752
rect 2504 -808 2548 -752
rect 4788 -760 4832 -752
rect 4900 -760 4920 -740
rect 4788 -800 4920 -760
rect 4788 -808 4832 -800
rect -180 -840 -60 -820
rect 4900 -820 4920 -800
rect 5000 -820 5020 -740
rect 4900 -840 5020 -820
rect -7588 -1155 -7516 -1142
rect -7588 -1289 -7575 -1155
rect -7529 -1289 -7516 -1155
rect -7588 -1302 -7516 -1289
rect -6386 -1155 -6314 -1142
rect -6386 -1289 -6373 -1155
rect -6327 -1289 -6314 -1155
rect -6386 -1302 -6314 -1289
rect -5600 -1180 -5480 -1160
rect -5600 -1260 -5580 -1180
rect -5500 -1200 -5480 -1180
rect 4900 -1180 5020 -1160
rect -5416 -1200 -5372 -1192
rect -5500 -1240 -5372 -1200
rect -5500 -1260 -5480 -1240
rect -5416 -1248 -5372 -1240
rect -892 -1248 -848 -1192
rect 264 -1248 308 -1192
rect 4788 -1200 4832 -1192
rect 4900 -1200 4920 -1180
rect 4788 -1240 4920 -1200
rect 4788 -1248 4832 -1240
rect -5600 -1280 -5480 -1260
rect 4900 -1260 4920 -1240
rect 5000 -1260 5020 -1180
rect 4900 -1280 5020 -1260
rect 5532 -1155 5604 -1142
rect 5532 -1289 5545 -1155
rect 5591 -1289 5604 -1155
rect 5532 -1302 5604 -1289
rect 6734 -1155 6806 -1142
rect 6734 -1289 6747 -1155
rect 6793 -1289 6806 -1155
rect 6734 -1302 6806 -1289
rect -6920 -2000 -6820 -1980
rect -6920 -2060 -6900 -2000
rect -6840 -2040 -6820 -2000
rect -6756 -2040 -6712 -2032
rect -6840 -2060 -6712 -2040
rect -6920 -2080 -6712 -2060
rect -6756 -2088 -6712 -2080
rect -3352 -2040 -3308 -2032
rect -3352 -2080 -3284 -2040
rect -3352 -2088 -3308 -2080
rect -6920 -2380 -6820 -2360
rect -6920 -2440 -6900 -2380
rect -6840 -2420 -6820 -2380
rect -6756 -2420 -6712 -2412
rect -6840 -2440 -6712 -2420
rect -6920 -2460 -6712 -2440
rect -6756 -2468 -6712 -2460
rect -3352 -2420 -3308 -2412
rect -3352 -2460 -3284 -2420
rect 6264 -2434 6320 -2390
rect -3352 -2468 -3308 -2460
rect 6264 -2654 6320 -2610
rect 6270 -2740 6310 -2654
rect 6210 -2760 6310 -2740
rect 6210 -2820 6230 -2760
rect 6290 -2820 6310 -2760
rect 6210 -2840 6310 -2820
rect 6210 -2920 6310 -2900
rect 6210 -2980 6230 -2920
rect 6290 -2980 6310 -2920
rect 6210 -3000 6310 -2980
rect 6270 -3052 6310 -3000
rect 6262 -3096 6318 -3052
rect -7204 -3473 -7004 -3460
rect -7204 -3519 -7191 -3473
rect -7017 -3519 -7004 -3473
rect -7204 -3582 -7004 -3519
rect -7204 -5145 -7004 -5082
rect -7204 -5191 -7191 -5145
rect -7017 -5191 -7004 -5145
rect -7204 -5204 -7004 -5191
rect -6344 -3473 -6144 -3460
rect -6344 -3519 -6331 -3473
rect -6157 -3519 -6144 -3473
rect -6344 -3582 -6144 -3519
rect -6344 -31645 -6144 -31582
rect -6344 -31691 -6331 -31645
rect -6157 -31691 -6144 -31645
rect -6344 -31704 -6144 -31691
rect -5544 -3473 -5344 -3460
rect -5544 -3519 -5531 -3473
rect -5357 -3519 -5344 -3473
rect -5544 -3582 -5344 -3519
rect -5544 -31645 -5344 -31582
rect -5544 -31691 -5531 -31645
rect -5357 -31691 -5344 -31645
rect -5544 -31704 -5344 -31691
rect -4744 -3473 -4544 -3460
rect -4744 -3519 -4731 -3473
rect -4557 -3519 -4544 -3473
rect -4744 -3582 -4544 -3519
rect -4744 -31645 -4544 -31582
rect -4744 -31691 -4731 -31645
rect -4557 -31691 -4544 -31645
rect -4744 -31704 -4544 -31691
rect -3944 -3473 -3744 -3460
rect -3944 -3519 -3931 -3473
rect -3757 -3519 -3744 -3473
rect -3944 -3582 -3744 -3519
rect -3944 -31645 -3744 -31582
rect -3944 -31691 -3931 -31645
rect -3757 -31691 -3744 -31645
rect -3944 -31704 -3744 -31691
rect -2344 -3473 -2144 -3460
rect -2344 -3519 -2331 -3473
rect -2157 -3519 -2144 -3473
rect -2344 -3582 -2144 -3519
rect -2344 -31645 -2144 -31582
rect -2344 -31691 -2331 -31645
rect -2157 -31691 -2144 -31645
rect -2344 -31704 -2144 -31691
rect -1544 -3473 -1344 -3460
rect -1544 -3519 -1531 -3473
rect -1357 -3519 -1344 -3473
rect -1544 -3582 -1344 -3519
rect -1544 -31645 -1344 -31582
rect -1544 -31691 -1531 -31645
rect -1357 -31691 -1344 -31645
rect -1544 -31704 -1344 -31691
rect 656 -3473 856 -3460
rect 656 -3519 669 -3473
rect 843 -3519 856 -3473
rect 656 -3582 856 -3519
rect 656 -31645 856 -31582
rect 656 -31691 669 -31645
rect 843 -31691 856 -31645
rect 656 -31704 856 -31691
rect 1456 -3473 1656 -3460
rect 1456 -3519 1469 -3473
rect 1643 -3519 1656 -3473
rect 1456 -3582 1656 -3519
rect 1456 -31645 1656 -31582
rect 1456 -31691 1469 -31645
rect 1643 -31691 1656 -31645
rect 1456 -31704 1656 -31691
rect 2256 -3473 2456 -3460
rect 2256 -3519 2269 -3473
rect 2443 -3519 2456 -3473
rect 2256 -3582 2456 -3519
rect 2256 -31645 2456 -31582
rect 2256 -31691 2269 -31645
rect 2443 -31691 2456 -31645
rect 2256 -31704 2456 -31691
rect 3056 -3473 3256 -3460
rect 3056 -3519 3069 -3473
rect 3243 -3519 3256 -3473
rect 3056 -3582 3256 -3519
rect 3056 -31645 3256 -31582
rect 3056 -31691 3069 -31645
rect 3243 -31691 3256 -31645
rect 3056 -31704 3256 -31691
rect 3856 -3473 4056 -3460
rect 3856 -3519 3869 -3473
rect 4043 -3519 4056 -3473
rect 3856 -3582 4056 -3519
rect 3856 -31645 4056 -31582
rect 3856 -31691 3869 -31645
rect 4043 -31691 4056 -31645
rect 3856 -31704 4056 -31691
rect 6262 -3316 6318 -3272
rect 5456 -3473 5656 -3460
rect 5456 -3519 5469 -3473
rect 5643 -3519 5656 -3473
rect 5456 -3582 5656 -3519
rect 5456 -31645 5656 -31582
rect 5456 -31691 5469 -31645
rect 5643 -31691 5656 -31645
rect 5456 -31704 5656 -31691
rect -6260 -31960 -6160 -31940
rect -6260 -32020 -6240 -31960
rect -6180 -32020 -6160 -31960
rect -6260 -32040 -6160 -32020
rect -5460 -31960 -5360 -31940
rect -5460 -32020 -5440 -31960
rect -5380 -32020 -5360 -31960
rect -5460 -32040 -5360 -32020
rect -4660 -31960 -4560 -31940
rect -4660 -32020 -4640 -31960
rect -4580 -32020 -4560 -31960
rect -4660 -32040 -4560 -32020
rect -3860 -31960 -3760 -31940
rect -3860 -32020 -3840 -31960
rect -3780 -32020 -3760 -31960
rect -3860 -32040 -3760 -32020
rect -2260 -31960 -2160 -31940
rect -2260 -32020 -2240 -31960
rect -2180 -32020 -2160 -31960
rect -2260 -32040 -2160 -32020
rect -1460 -31960 -1360 -31940
rect -1460 -32020 -1440 -31960
rect -1380 -32020 -1360 -31960
rect -1460 -32040 -1360 -32020
rect 680 -31960 780 -31940
rect 680 -32020 700 -31960
rect 760 -32020 780 -31960
rect 680 -32040 780 -32020
rect 1480 -31960 1580 -31940
rect 1480 -32020 1500 -31960
rect 1560 -32020 1580 -31960
rect 1480 -32040 1580 -32020
rect 2280 -31960 2380 -31940
rect 2280 -32020 2300 -31960
rect 2360 -32020 2380 -31960
rect 2280 -32040 2380 -32020
rect 3080 -31960 3180 -31940
rect 3080 -32020 3100 -31960
rect 3160 -32020 3180 -31960
rect 3080 -32040 3180 -32020
rect 3880 -31960 3980 -31940
rect 3880 -32020 3900 -31960
rect 3960 -32020 3980 -31960
rect 3880 -32040 3980 -32020
rect 5480 -31960 5580 -31940
rect 5480 -32020 5500 -31960
rect 5560 -32020 5580 -31960
rect 5480 -32040 5580 -32020
rect -6260 -32104 -6220 -32040
rect -5460 -32104 -5420 -32040
rect -4660 -32104 -4620 -32040
rect -3860 -32104 -3820 -32040
rect -2260 -32100 -2220 -32040
rect -1460 -32100 -1420 -32040
rect -6268 -32148 -6212 -32104
rect -5468 -32148 -5412 -32104
rect -4668 -32148 -4612 -32104
rect -3868 -32148 -3812 -32104
rect -2268 -32144 -2212 -32100
rect -1468 -32144 -1412 -32100
rect 740 -32108 780 -32040
rect 1540 -32108 1580 -32040
rect 2340 -32108 2380 -32040
rect 3140 -32108 3180 -32040
rect 3940 -32108 3980 -32040
rect 5540 -32100 5580 -32040
rect -6268 -32976 -6212 -32932
rect -5468 -32976 -5412 -32932
rect -4668 -32976 -4612 -32932
rect -3868 -32976 -3812 -32932
rect 732 -32152 788 -32108
rect 1532 -32152 1588 -32108
rect 2332 -32152 2388 -32108
rect 3132 -32152 3188 -32108
rect 3932 -32152 3988 -32108
rect 5532 -32144 5588 -32100
rect 5532 -32356 5588 -32312
rect 732 -32756 788 -32712
rect 1532 -32756 1588 -32712
rect 2332 -32756 2388 -32712
rect 3132 -32756 3188 -32712
rect 3932 -32756 3988 -32712
rect -2268 -33756 -2212 -33712
rect -1468 -33756 -1412 -33712
rect -6344 -34173 -6144 -34160
rect -6344 -34219 -6331 -34173
rect -6157 -34219 -6144 -34173
rect -6344 -34282 -6144 -34219
rect -6344 -62345 -6144 -62282
rect -6344 -62391 -6331 -62345
rect -6157 -62391 -6144 -62345
rect -6344 -62404 -6144 -62391
rect -5544 -34173 -5344 -34160
rect -5544 -34219 -5531 -34173
rect -5357 -34219 -5344 -34173
rect -5544 -34282 -5344 -34219
rect -5544 -62345 -5344 -62282
rect -5544 -62391 -5531 -62345
rect -5357 -62391 -5344 -62345
rect -5544 -62404 -5344 -62391
rect -4744 -34173 -4544 -34160
rect -4744 -34219 -4731 -34173
rect -4557 -34219 -4544 -34173
rect -4744 -34282 -4544 -34219
rect -4744 -62345 -4544 -62282
rect -4744 -62391 -4731 -62345
rect -4557 -62391 -4544 -62345
rect -4744 -62404 -4544 -62391
rect -3944 -34173 -3744 -34160
rect -3944 -34219 -3931 -34173
rect -3757 -34219 -3744 -34173
rect -3944 -34282 -3744 -34219
rect -3944 -62345 -3744 -62282
rect -3944 -62391 -3931 -62345
rect -3757 -62391 -3744 -62345
rect -3944 -62404 -3744 -62391
rect -2344 -34180 -2260 -34160
rect -2160 -34180 -2144 -34160
rect -2344 -34282 -2144 -34180
rect -2344 -62345 -2144 -62282
rect -2344 -62391 -2331 -62345
rect -2157 -62391 -2144 -62345
rect -2344 -62404 -2144 -62391
rect -1544 -34173 -1344 -34160
rect -1544 -34219 -1531 -34173
rect -1357 -34219 -1344 -34173
rect -1544 -34282 -1344 -34219
rect -1544 -62345 -1344 -62282
rect -1544 -62391 -1531 -62345
rect -1357 -62391 -1344 -62345
rect -1544 -62404 -1344 -62391
rect 656 -34133 856 -34120
rect 656 -34179 669 -34133
rect 843 -34179 856 -34133
rect 656 -34242 856 -34179
rect 656 -62305 856 -62242
rect 656 -62351 669 -62305
rect 843 -62351 856 -62305
rect 656 -62364 856 -62351
rect 1456 -34133 1656 -34120
rect 1456 -34179 1469 -34133
rect 1643 -34179 1656 -34133
rect 1456 -34242 1656 -34179
rect 1456 -62305 1656 -62242
rect 1456 -62351 1469 -62305
rect 1643 -62351 1656 -62305
rect 1456 -62364 1656 -62351
rect 2256 -34133 2456 -34120
rect 2256 -34179 2269 -34133
rect 2443 -34179 2456 -34133
rect 2256 -34242 2456 -34179
rect 2256 -62305 2456 -62242
rect 2256 -62351 2269 -62305
rect 2443 -62351 2456 -62305
rect 2256 -62364 2456 -62351
rect 3056 -34133 3256 -34120
rect 3056 -34179 3069 -34133
rect 3243 -34179 3256 -34133
rect 3056 -34242 3256 -34179
rect 3056 -62305 3256 -62242
rect 3056 -62351 3069 -62305
rect 3243 -62351 3256 -62305
rect 3056 -62364 3256 -62351
rect 3856 -34133 4056 -34120
rect 3856 -34179 3869 -34133
rect 4043 -34179 4056 -34133
rect 3856 -34242 4056 -34179
rect 3856 -62305 4056 -62242
rect 3856 -62351 3869 -62305
rect 4043 -62351 4056 -62305
rect 3856 -62364 4056 -62351
rect 5456 -34133 5656 -34120
rect 5456 -34179 5469 -34133
rect 5643 -34179 5656 -34133
rect 5456 -34242 5656 -34179
rect 5456 -62305 5656 -62242
rect 5456 -62351 5469 -62305
rect 5643 -62351 5656 -62305
rect 5456 -62364 5656 -62351
<< polycontact >>
rect -5580 -820 -5500 -740
rect -520 -820 -440 -740
rect -160 -820 -80 -740
rect 4920 -820 5000 -740
rect -7575 -1289 -7529 -1155
rect -6373 -1289 -6327 -1155
rect -5580 -1260 -5500 -1180
rect 4920 -1260 5000 -1180
rect 5545 -1289 5591 -1155
rect 6747 -1289 6793 -1155
rect -6900 -2060 -6840 -2000
rect -6900 -2440 -6840 -2380
rect 6230 -2820 6290 -2760
rect 6230 -2980 6290 -2920
rect -7191 -3519 -7017 -3473
rect -7191 -5191 -7017 -5145
rect -6331 -3519 -6157 -3473
rect -6331 -31691 -6157 -31645
rect -5531 -3519 -5357 -3473
rect -5531 -31691 -5357 -31645
rect -4731 -3519 -4557 -3473
rect -4731 -31691 -4557 -31645
rect -3931 -3519 -3757 -3473
rect -3931 -31691 -3757 -31645
rect -2331 -3519 -2157 -3473
rect -2331 -31691 -2157 -31645
rect -1531 -3519 -1357 -3473
rect -1531 -31691 -1357 -31645
rect 669 -3519 843 -3473
rect 669 -31691 843 -31645
rect 1469 -3519 1643 -3473
rect 1469 -31691 1643 -31645
rect 2269 -3519 2443 -3473
rect 2269 -31691 2443 -31645
rect 3069 -3519 3243 -3473
rect 3069 -31691 3243 -31645
rect 3869 -3519 4043 -3473
rect 3869 -31691 4043 -31645
rect 5469 -3519 5643 -3473
rect 5469 -31691 5643 -31645
rect -6240 -32020 -6180 -31960
rect -5440 -32020 -5380 -31960
rect -4640 -32020 -4580 -31960
rect -3840 -32020 -3780 -31960
rect -2240 -32020 -2180 -31960
rect -1440 -32020 -1380 -31960
rect 700 -32020 760 -31960
rect 1500 -32020 1560 -31960
rect 2300 -32020 2360 -31960
rect 3100 -32020 3160 -31960
rect 3900 -32020 3960 -31960
rect 5500 -32020 5560 -31960
rect -6331 -34219 -6157 -34173
rect -6331 -62391 -6157 -62345
rect -5531 -34219 -5357 -34173
rect -5531 -62391 -5357 -62345
rect -4731 -34219 -4557 -34173
rect -4731 -62391 -4557 -62345
rect -3931 -34219 -3757 -34173
rect -3931 -62391 -3757 -62345
rect -2331 -62391 -2157 -62345
rect -1531 -34219 -1357 -34173
rect -1531 -62391 -1357 -62345
rect 669 -34179 843 -34133
rect 669 -62351 843 -62305
rect 1469 -34179 1643 -34133
rect 1469 -62351 1643 -62305
rect 2269 -34179 2443 -34133
rect 2269 -62351 2443 -62305
rect 3069 -34179 3243 -34133
rect 3069 -62351 3243 -62305
rect 3869 -34179 4043 -34133
rect 3869 -62351 4043 -62305
rect 5469 -34179 5643 -34133
rect 5469 -62351 5643 -62305
<< ppolysilicide >>
rect -7516 -1302 -6386 -1142
rect 5604 -1302 6734 -1142
<< nhighres >>
rect -7204 -5082 -7004 -3582
rect -6344 -31582 -6144 -3582
rect -5544 -31582 -5344 -3582
rect -4744 -31582 -4544 -3582
rect -3944 -31582 -3744 -3582
rect -2344 -31582 -2144 -3582
rect -1544 -31582 -1344 -3582
rect 656 -31582 856 -3582
rect 1456 -31582 1656 -3582
rect 2256 -31582 2456 -3582
rect 3056 -31582 3256 -3582
rect 3856 -31582 4056 -3582
rect 5456 -31582 5656 -3582
rect -6344 -62282 -6144 -34282
rect -5544 -62282 -5344 -34282
rect -4744 -62282 -4544 -34282
rect -3944 -62282 -3744 -34282
rect -2344 -62282 -2144 -34282
rect -1544 -62282 -1344 -34282
rect 656 -62242 856 -34242
rect 1456 -62242 1656 -34242
rect 2256 -62242 2456 -34242
rect 3056 -62242 3256 -34242
rect 3856 -62242 4056 -34242
rect 5456 -62242 5656 -34242
<< pdiffres >>
rect -1768 66 -848 266
rect 252 66 1172 266
<< metal1 >>
rect -380 1060 -220 1520
rect -380 960 -350 1060
rect -250 960 -220 1060
rect -1881 253 -1835 264
rect -3220 80 -1881 240
rect -3220 -380 -3140 80
rect -1881 68 -1835 79
rect -781 253 -735 264
rect -380 240 -220 960
rect 5100 780 5220 800
rect 5100 700 5120 780
rect 5200 700 5220 780
rect 139 253 185 264
rect -735 80 139 240
rect -781 68 -735 79
rect 139 68 185 79
rect 1239 253 1285 264
rect 1285 80 2640 240
rect 1239 68 1285 79
rect -8260 -400 -3140 -380
rect 2560 -220 2640 80
rect 2620 -300 2640 -220
rect -8260 -480 140 -400
rect -8260 -500 -3140 -480
rect -5360 -677 -5280 -660
rect -3220 -677 -3140 -500
rect -760 -560 -640 -540
rect -760 -620 -740 -560
rect -660 -620 -640 -560
rect -760 -677 -640 -620
rect -6360 -740 -5500 -720
rect -5370 -723 -5359 -677
rect -3145 -723 -3134 -677
rect -2910 -723 -2899 -677
rect -685 -720 -640 -677
rect -360 -560 -240 -540
rect -360 -620 -340 -560
rect -260 -620 -240 -560
rect -685 -723 -674 -720
rect -360 -740 -240 -620
rect 60 -677 140 -480
rect 2560 -677 2640 -300
rect 50 -723 61 -677
rect 2275 -723 2286 -677
rect 2550 -723 2561 -677
rect 4775 -723 4786 -677
rect 5100 -720 5220 700
rect 4920 -740 7340 -720
rect -6360 -820 -6340 -740
rect -6260 -820 -5580 -740
rect -540 -820 -520 -740
rect -440 -820 -160 -740
rect -80 -820 -60 -740
rect 5000 -820 7340 -740
rect -6360 -840 -5500 -820
rect -5440 -883 -5359 -837
rect -3145 -883 -2899 -837
rect -685 -883 -674 -837
rect 50 -883 61 -837
rect 2275 -883 2561 -837
rect 4775 -883 4860 -837
rect 4920 -840 7340 -820
rect -5440 -1117 -5370 -883
rect -5320 -980 -5300 -934
rect -3160 -980 -2884 -934
rect -744 -940 -724 -934
rect -744 -980 -700 -940
rect 100 -980 120 -934
rect 2260 -980 2576 -934
rect 4716 -980 4736 -934
rect -800 -1020 -700 -980
rect -800 -1080 -780 -1020
rect -720 -1080 -700 -1020
rect 80 -1020 180 -980
rect 80 -1080 100 -1020
rect 160 -1080 180 -1020
rect 4800 -1117 4860 -883
rect -7575 -1155 -7529 -1144
rect -8260 -1280 -7575 -1160
rect -7575 -1300 -7529 -1289
rect -6373 -1155 -6327 -1144
rect -6327 -1180 -5500 -1160
rect -5440 -1163 -5359 -1117
rect -905 -1163 -894 -1117
rect 310 -1163 321 -1117
rect 4775 -1163 4860 -1117
rect 5545 -1155 5591 -1144
rect -6327 -1260 -5580 -1180
rect -6327 -1280 -5500 -1260
rect 4920 -1180 5545 -1160
rect 5000 -1260 5545 -1180
rect -6373 -1300 -6327 -1289
rect -5780 -1540 -5680 -1280
rect -5370 -1323 -5359 -1277
rect -905 -1323 321 -1277
rect 4775 -1323 4786 -1277
rect 4920 -1280 5545 -1260
rect -5320 -1420 -5300 -1374
rect -905 -1380 -894 -1374
rect -905 -1420 -780 -1380
rect -940 -1440 -780 -1420
rect -720 -1440 -700 -1380
rect -940 -1460 -700 -1440
rect -5780 -1580 -2060 -1540
rect -5780 -1640 -2140 -1580
rect -2080 -1640 -2060 -1580
rect -940 -1600 -820 -1580
rect -940 -1660 -920 -1600
rect -840 -1660 -820 -1600
rect -6700 -1880 -2960 -1800
rect -6700 -1957 -3360 -1880
rect -6920 -2000 -6820 -1980
rect -6920 -2060 -6900 -2000
rect -6840 -2060 -6820 -2000
rect -6710 -2003 -6699 -1957
rect -3365 -2003 -3354 -1957
rect -6920 -2180 -6820 -2060
rect -6710 -2163 -6699 -2117
rect -3365 -2140 -3354 -2117
rect -3365 -2163 -3360 -2160
rect -7180 -2260 -6820 -2180
rect -7180 -2620 -7020 -2260
rect -6920 -2380 -6820 -2260
rect -6700 -2220 -3360 -2163
rect -3260 -2220 -3180 -2200
rect -6700 -2227 -3240 -2220
rect -6700 -2273 -6660 -2227
rect -3380 -2273 -3240 -2227
rect -6700 -2280 -3240 -2273
rect -6700 -2337 -3360 -2280
rect -3260 -2300 -3180 -2280
rect -6920 -2440 -6900 -2380
rect -6840 -2440 -6820 -2380
rect -6710 -2383 -6699 -2337
rect -3365 -2383 -3354 -2337
rect -6920 -2460 -6820 -2440
rect -6710 -2543 -6699 -2497
rect -3365 -2520 -3354 -2497
rect -3365 -2543 -3284 -2520
rect -6640 -2620 -6480 -2543
rect -3400 -2580 -3284 -2543
rect -7180 -2700 -6480 -2620
rect -7180 -3473 -7020 -2700
rect -5080 -3120 -5000 -3100
rect -5080 -3180 -5060 -3120
rect -5080 -3460 -5000 -3180
rect -6340 -3473 -3740 -3460
rect -7202 -3519 -7191 -3473
rect -7017 -3519 -7006 -3473
rect -6342 -3519 -6331 -3473
rect -6157 -3519 -5531 -3473
rect -5357 -3519 -4731 -3473
rect -4557 -3519 -3931 -3473
rect -3757 -3519 -3740 -3473
rect -7180 -3520 -7020 -3519
rect -6340 -3520 -3740 -3519
rect -7202 -5191 -7191 -5145
rect -7017 -5191 -7006 -5145
rect -7180 -6160 -7020 -5191
rect -7180 -6280 -7160 -6160
rect -7040 -6280 -7020 -6160
rect -7180 -62680 -7020 -6280
rect -6260 -31645 -6160 -31640
rect -5460 -31645 -5360 -31640
rect -4660 -31645 -4560 -31640
rect -3860 -31645 -3760 -31640
rect -6342 -31691 -6331 -31645
rect -6157 -31691 -6146 -31645
rect -5542 -31691 -5531 -31645
rect -5357 -31691 -5346 -31645
rect -4742 -31691 -4731 -31645
rect -4557 -31691 -4546 -31645
rect -3942 -31691 -3931 -31645
rect -3757 -31691 -3746 -31645
rect -6260 -31960 -6160 -31691
rect -6260 -32020 -6240 -31960
rect -6180 -32020 -6160 -31960
rect -6260 -32040 -6160 -32020
rect -5460 -31960 -5360 -31691
rect -5460 -32020 -5440 -31960
rect -5380 -32020 -5360 -31960
rect -5460 -32040 -5360 -32020
rect -4660 -31960 -4560 -31691
rect -4660 -32020 -4640 -31960
rect -4580 -32020 -4560 -31960
rect -4660 -32040 -4560 -32020
rect -3860 -31960 -3760 -31691
rect -3860 -32020 -3840 -31960
rect -3780 -32020 -3760 -31960
rect -3860 -32040 -3760 -32020
rect -3120 -32100 -2960 -1880
rect -940 -1960 -820 -1660
rect -940 -2020 -920 -1960
rect -840 -2020 -820 -1960
rect -940 -2080 -820 -2020
rect -380 -2080 -220 -1323
rect 310 -1380 321 -1374
rect 80 -1440 100 -1380
rect 160 -1420 321 -1380
rect 4716 -1420 4736 -1374
rect 160 -1440 360 -1420
rect 80 -1460 360 -1440
rect 1460 -1560 4160 -1540
rect 1460 -1580 4100 -1560
rect 220 -1600 340 -1580
rect 220 -1660 240 -1600
rect 320 -1660 340 -1600
rect 1460 -1640 1480 -1580
rect 1540 -1620 4100 -1580
rect 1540 -1640 4160 -1620
rect 220 -1960 340 -1660
rect 220 -2020 240 -1960
rect 320 -2020 340 -1960
rect 220 -2080 340 -2020
rect -940 -2180 340 -2080
rect -2840 -2220 -2740 -2200
rect -2840 -2280 -2820 -2220
rect -2760 -2280 -2740 -2220
rect -2840 -2300 -2740 -2280
rect -940 -2300 -820 -2180
rect -2820 -2800 -2760 -2300
rect -940 -2360 -920 -2300
rect -840 -2360 -820 -2300
rect -940 -2660 -820 -2360
rect -940 -2720 -920 -2660
rect -840 -2720 -820 -2660
rect -940 -2740 -820 -2720
rect -700 -2780 -600 -2760
rect -700 -2800 -680 -2780
rect -2820 -2840 -680 -2800
rect -620 -2840 -600 -2780
rect -2820 -2860 -600 -2840
rect -1880 -2940 -1800 -2920
rect -1880 -3000 -1860 -2940
rect -1880 -3460 -1800 -3000
rect -2340 -3473 -1340 -3460
rect -2342 -3519 -2331 -3473
rect -2157 -3519 -1531 -3473
rect -1357 -3519 -1340 -3473
rect -2340 -3520 -1340 -3519
rect -2260 -31645 -2160 -31640
rect -1460 -31645 -1360 -31640
rect -2342 -31691 -2331 -31645
rect -2157 -31691 -2146 -31645
rect -1542 -31691 -1531 -31645
rect -1357 -31691 -1346 -31645
rect -2260 -31960 -2160 -31691
rect -2260 -32020 -2240 -31960
rect -2180 -32020 -2160 -31960
rect -2260 -32040 -2160 -32020
rect -1460 -31960 -1360 -31691
rect -1460 -32020 -1440 -31960
rect -1380 -32020 -1360 -31960
rect -1460 -32040 -1360 -32020
rect -6860 -32160 -6297 -32100
rect -6860 -34480 -6700 -32160
rect -6343 -32161 -6297 -32160
rect -6440 -32220 -6394 -32206
rect -6440 -32980 -6394 -32919
rect -6343 -32930 -6297 -32919
rect -6183 -32160 -5497 -32100
rect -6183 -32161 -6137 -32160
rect -5543 -32161 -5497 -32160
rect -6183 -32930 -6137 -32919
rect -5640 -32220 -5594 -32206
rect -5640 -32980 -5594 -32919
rect -5543 -32930 -5497 -32919
rect -5383 -32160 -4697 -32100
rect -5383 -32161 -5337 -32160
rect -4743 -32161 -4697 -32160
rect -5383 -32930 -5337 -32919
rect -4840 -32220 -4794 -32206
rect -4840 -32980 -4794 -32919
rect -4743 -32930 -4697 -32919
rect -4583 -32160 -3897 -32100
rect -4583 -32161 -4537 -32160
rect -3943 -32161 -3897 -32160
rect -4583 -32930 -4537 -32919
rect -4040 -32220 -3994 -32206
rect -4040 -32980 -3994 -32919
rect -3943 -32930 -3897 -32919
rect -3783 -32146 -2297 -32100
rect -3783 -32160 -2480 -32146
rect -2343 -32157 -2297 -32146
rect -3783 -32161 -3737 -32160
rect -3783 -32930 -3737 -32919
rect -2446 -32220 -2400 -32200
rect -6440 -33820 -6380 -32980
rect -5640 -33820 -5580 -32980
rect -4840 -33820 -4780 -32980
rect -4040 -33820 -3980 -32980
rect -2446 -33820 -2400 -33699
rect -2343 -33710 -2297 -33699
rect -2183 -32146 -1497 -32092
rect -380 -32140 -220 -2180
rect 220 -2300 340 -2180
rect 220 -2360 240 -2300
rect 320 -2360 340 -2300
rect 220 -2660 340 -2360
rect 220 -2720 240 -2660
rect 320 -2720 340 -2660
rect 220 -2740 340 -2720
rect -100 -2780 0 -2760
rect -100 -2840 -80 -2780
rect -20 -2800 0 -2780
rect 4420 -2800 4520 -1420
rect 5080 -1540 5180 -1280
rect 5545 -1300 5591 -1289
rect 6747 -1155 6793 -1144
rect 6793 -1280 7340 -1160
rect 6747 -1300 6793 -1289
rect 4780 -1560 5180 -1540
rect 4840 -1620 5180 -1560
rect 4780 -1640 5180 -1620
rect -20 -2840 4520 -2800
rect -100 -2860 4520 -2840
rect 2320 -3120 2400 -3100
rect 2320 -3180 2340 -3120
rect 2320 -3460 2400 -3180
rect 660 -3473 4060 -3460
rect 660 -3519 669 -3473
rect 843 -3519 1469 -3473
rect 1643 -3519 2269 -3473
rect 2443 -3519 3069 -3473
rect 3243 -3519 3869 -3473
rect 4043 -3519 4060 -3473
rect 660 -3520 4060 -3519
rect 4420 -3960 4520 -2860
rect 4420 -4020 4460 -3960
rect 4420 -4040 4520 -4020
rect 4700 -1940 7340 -1780
rect 680 -31645 780 -31640
rect 1480 -31645 1580 -31640
rect 2280 -31645 2380 -31640
rect 3080 -31645 3180 -31640
rect 3880 -31645 3980 -31640
rect 658 -31691 669 -31645
rect 843 -31691 854 -31645
rect 1458 -31691 1469 -31645
rect 1643 -31691 1654 -31645
rect 2258 -31691 2269 -31645
rect 2443 -31691 2454 -31645
rect 3058 -31691 3069 -31645
rect 3243 -31691 3254 -31645
rect 3858 -31691 3869 -31645
rect 4043 -31691 4054 -31645
rect 680 -31960 780 -31691
rect 680 -32020 700 -31960
rect 760 -32020 780 -31960
rect 680 -32040 780 -32020
rect 1480 -31960 1580 -31691
rect 1480 -32020 1500 -31960
rect 1560 -32020 1580 -31960
rect 1480 -32040 1580 -32020
rect 2280 -31960 2380 -31691
rect 2280 -32020 2300 -31960
rect 2360 -32020 2380 -31960
rect 2280 -32040 2380 -32020
rect 3080 -31960 3180 -31691
rect 3080 -32020 3100 -31960
rect 3160 -32020 3180 -31960
rect 3080 -32040 3180 -32020
rect 3880 -31960 3980 -31691
rect 3880 -32020 3900 -31960
rect 3960 -32020 3980 -31960
rect 3880 -32040 3980 -32020
rect 4700 -32100 4860 -1940
rect 6085 -2220 6250 -2200
rect 6085 -2280 6170 -2220
rect 6230 -2280 6250 -2220
rect 6085 -2300 6250 -2280
rect 6085 -2436 6150 -2300
rect 6085 -2447 6235 -2436
rect 6131 -2597 6189 -2447
rect 6085 -2608 6235 -2597
rect 6349 -2440 6395 -2436
rect 6349 -2447 6410 -2440
rect 6395 -2597 6410 -2447
rect 6349 -2608 6410 -2597
rect 6350 -2640 6410 -2608
rect 6350 -2680 6430 -2640
rect 6210 -2760 6310 -2740
rect 6210 -2820 6230 -2760
rect 6290 -2820 6310 -2760
rect 5500 -2840 5600 -2820
rect 6210 -2840 6310 -2820
rect 5500 -2900 5520 -2840
rect 5580 -2900 6310 -2840
rect 5500 -2920 5600 -2900
rect 5520 -3473 5600 -2920
rect 6210 -2920 6310 -2900
rect 6210 -2980 6230 -2920
rect 6290 -2980 6310 -2920
rect 6210 -3000 6310 -2980
rect 6370 -2820 6430 -2680
rect 6370 -2840 6570 -2820
rect 6370 -2900 6490 -2840
rect 6550 -2900 6570 -2840
rect 6370 -2920 6570 -2900
rect 6370 -3080 6430 -2920
rect 6350 -3098 6430 -3080
rect 6080 -3109 6233 -3098
rect 6080 -3259 6084 -3109
rect 6130 -3259 6187 -3109
rect 6080 -3270 6233 -3259
rect 6347 -3109 6430 -3098
rect 6393 -3120 6430 -3109
rect 6393 -3259 6410 -3120
rect 6347 -3260 6410 -3259
rect 6347 -3270 6393 -3260
rect 5458 -3519 5469 -3473
rect 5643 -3519 5654 -3473
rect 5520 -3520 5600 -3519
rect 6080 -3620 6180 -3270
rect 6080 -3940 6220 -3620
rect 6080 -3960 7420 -3940
rect 6080 -4020 6120 -3960
rect 6180 -4020 7420 -3960
rect 6080 -4040 7420 -4020
rect 5480 -31645 5580 -31640
rect 5458 -31691 5469 -31645
rect 5643 -31691 5654 -31645
rect 5480 -31960 5580 -31691
rect 5480 -32020 5500 -31960
rect 5560 -32020 5580 -31960
rect 5480 -32040 5580 -32020
rect -1380 -32146 -220 -32140
rect -2183 -32157 -2137 -32146
rect -1543 -32157 -1497 -32146
rect -2183 -33710 -2137 -33699
rect -1646 -32220 -1600 -32200
rect -1646 -33820 -1600 -33699
rect -1543 -33710 -1497 -33699
rect -1383 -32157 -220 -32146
rect 817 -32154 1503 -32100
rect 1617 -32154 2303 -32100
rect 2417 -32154 3103 -32100
rect 3217 -32154 3903 -32100
rect -1337 -32160 -220 -32157
rect -1337 -32680 657 -32160
rect 3057 -32165 3103 -32160
rect -1337 -33699 -1300 -32680
rect 620 -32699 657 -32680
rect 620 -32700 703 -32699
rect 657 -32710 703 -32700
rect 863 -32220 966 -32200
rect 863 -32699 920 -32220
rect 817 -32710 966 -32699
rect 1457 -32710 1503 -32699
rect 1663 -32220 1766 -32200
rect 1663 -32699 1720 -32220
rect 1617 -32710 1766 -32699
rect 2257 -32710 2303 -32699
rect 2463 -32220 2566 -32200
rect 2463 -32699 2520 -32220
rect 2417 -32710 2566 -32699
rect 3057 -32710 3103 -32699
rect 3217 -32165 3263 -32154
rect 3900 -32165 3903 -32154
rect 3263 -32220 3366 -32200
rect 3263 -32699 3320 -32220
rect 3217 -32710 3366 -32699
rect 3857 -32710 3903 -32699
rect 4017 -32152 5503 -32100
rect 4017 -32165 4063 -32152
rect 5457 -32157 5503 -32152
rect 4063 -32220 4166 -32200
rect 4063 -32699 4120 -32220
rect 5457 -32310 5503 -32299
rect 5617 -32152 6340 -32100
rect 5617 -32157 5663 -32152
rect 5663 -32211 5766 -32200
rect 5663 -32299 5720 -32211
rect 5617 -32310 5766 -32299
rect 4017 -32710 4166 -32699
rect -1383 -33700 -1300 -33699
rect 920 -32760 966 -32710
rect 1720 -32760 1766 -32710
rect 2520 -32760 2566 -32710
rect 3320 -32760 3366 -32710
rect 4120 -32760 4166 -32710
rect 5720 -32360 5766 -32310
rect -1383 -33710 -1337 -33700
rect 920 -33780 980 -32760
rect 1720 -33780 1780 -32760
rect 2520 -33780 2580 -32760
rect 3320 -33780 3380 -32760
rect 4120 -33780 4180 -32760
rect 5720 -33780 5780 -32360
rect -6440 -33880 -6200 -33820
rect -5640 -33880 -5400 -33820
rect -4840 -33880 -4600 -33820
rect -4040 -33880 -3800 -33820
rect -2446 -33880 -2200 -33820
rect -1646 -33880 -1400 -33820
rect -6280 -34160 -6200 -33880
rect -5480 -34160 -5400 -33880
rect -4680 -34160 -4600 -33880
rect -3880 -34160 -3800 -33880
rect -6280 -34173 -6160 -34160
rect -5480 -34173 -5360 -34160
rect -4680 -34173 -4560 -34160
rect -3880 -34173 -3760 -34160
rect -2280 -34173 -2200 -33880
rect -1480 -34160 -1400 -33880
rect 720 -33860 980 -33780
rect 1520 -33860 1780 -33780
rect 2320 -33860 2580 -33780
rect 3120 -33860 3380 -33780
rect 3920 -33860 4180 -33780
rect 5520 -33860 5780 -33780
rect 6180 -33340 6340 -32152
rect 6900 -33340 7000 -4040
rect 6180 -33500 7000 -33340
rect 720 -34120 800 -33860
rect 1520 -34120 1600 -33860
rect 2320 -34120 2400 -33860
rect 3120 -34120 3200 -33860
rect 3920 -34120 4000 -33860
rect 5520 -34120 5600 -33860
rect 720 -34133 840 -34120
rect 1520 -34133 1640 -34120
rect 2320 -34133 2440 -34120
rect 3120 -34133 3240 -34120
rect 3920 -34133 4040 -34120
rect 5520 -34133 5640 -34120
rect -1480 -34173 -1360 -34160
rect -6342 -34219 -6331 -34173
rect -6157 -34219 -6146 -34173
rect -5542 -34219 -5531 -34173
rect -5357 -34219 -5346 -34173
rect -4742 -34219 -4731 -34173
rect -4557 -34219 -4546 -34173
rect -3942 -34219 -3931 -34173
rect -3757 -34219 -3746 -34173
rect -6260 -34220 -6160 -34219
rect -5460 -34220 -5360 -34219
rect -4660 -34220 -4560 -34219
rect -3860 -34220 -3760 -34219
rect -2260 -34220 -2160 -34180
rect -1542 -34219 -1531 -34173
rect -1357 -34219 -1346 -34173
rect 658 -34179 669 -34133
rect 843 -34179 854 -34133
rect 1458 -34179 1469 -34133
rect 1643 -34179 1654 -34133
rect 2258 -34179 2269 -34133
rect 2443 -34179 2454 -34133
rect 3058 -34179 3069 -34133
rect 3243 -34179 3254 -34133
rect 3858 -34179 3869 -34133
rect 4043 -34179 4054 -34133
rect 5458 -34179 5469 -34133
rect 5643 -34179 5654 -34133
rect 740 -34180 840 -34179
rect 1540 -34180 1640 -34179
rect 2340 -34180 2440 -34179
rect 3140 -34180 3240 -34179
rect 3940 -34180 4040 -34179
rect 5540 -34180 5640 -34179
rect -1460 -34220 -1360 -34219
rect 6180 -34480 6340 -33500
rect -6860 -34640 6340 -34480
rect 740 -62305 840 -62300
rect 1540 -62305 1640 -62300
rect 2340 -62305 2440 -62300
rect 3140 -62305 3240 -62300
rect 3940 -62305 4040 -62300
rect 5540 -62305 5640 -62300
rect -6260 -62345 -6160 -62340
rect -5460 -62345 -5360 -62340
rect -4660 -62345 -4560 -62340
rect -3860 -62345 -3760 -62340
rect -2260 -62345 -2160 -62340
rect -1460 -62345 -1360 -62340
rect -6342 -62391 -6331 -62345
rect -6157 -62391 -6146 -62345
rect -5542 -62391 -5531 -62345
rect -5357 -62391 -5346 -62345
rect -4742 -62391 -4731 -62345
rect -4557 -62391 -4546 -62345
rect -3942 -62391 -3931 -62345
rect -3757 -62391 -3746 -62345
rect -2342 -62391 -2331 -62345
rect -2157 -62391 -2146 -62345
rect -1542 -62391 -1531 -62345
rect -1357 -62391 -1346 -62345
rect 658 -62351 669 -62305
rect 843 -62351 854 -62305
rect 1458 -62351 1469 -62305
rect 1643 -62351 1654 -62305
rect 2258 -62351 2269 -62305
rect 2443 -62351 2454 -62305
rect 3058 -62351 3069 -62305
rect 3243 -62351 3254 -62305
rect 3858 -62351 3869 -62305
rect 4043 -62351 4054 -62305
rect 5458 -62351 5469 -62305
rect 5643 -62351 5654 -62305
rect -6260 -62680 -6160 -62391
rect -5460 -62680 -5360 -62391
rect -4660 -62680 -4560 -62391
rect -3860 -62680 -3760 -62391
rect -2260 -62680 -2160 -62391
rect -1460 -62680 -1360 -62391
rect 740 -62680 840 -62351
rect 1540 -62680 1640 -62351
rect 2340 -62680 2440 -62351
rect 3140 -62680 3240 -62351
rect 3940 -62680 4040 -62351
rect 5540 -62680 5640 -62351
rect -7180 -62720 6660 -62680
rect -7180 -62800 6540 -62720
rect 6620 -62800 6660 -62720
rect -7180 -62840 6660 -62800
<< via1 >>
rect -350 960 -250 1060
rect 5120 700 5200 780
rect 2560 -300 2620 -220
rect -740 -620 -660 -560
rect -340 -620 -260 -560
rect -6340 -820 -6260 -740
rect -780 -1080 -720 -1020
rect 100 -1080 160 -1020
rect -780 -1440 -720 -1380
rect -2140 -1640 -2080 -1580
rect -920 -1660 -840 -1600
rect -3240 -2280 -3180 -2220
rect -5060 -3180 -5000 -3120
rect -7160 -6280 -7040 -6160
rect -920 -2020 -840 -1960
rect 100 -1440 160 -1380
rect 240 -1660 320 -1600
rect 1480 -1640 1540 -1580
rect 4100 -1620 4160 -1560
rect 240 -2020 320 -1960
rect -2820 -2280 -2760 -2220
rect -920 -2360 -840 -2300
rect -920 -2720 -840 -2660
rect -680 -2840 -620 -2780
rect -1860 -3000 -1800 -2940
rect 240 -2360 320 -2300
rect 240 -2720 320 -2660
rect -80 -2840 -20 -2780
rect 4780 -1620 4840 -1560
rect 2340 -3180 2400 -3120
rect 4460 -4020 4520 -3960
rect 6170 -2280 6230 -2220
rect 5520 -2900 5580 -2840
rect 6490 -2900 6550 -2840
rect 6120 -4020 6180 -3960
rect 6540 -62800 6620 -62720
<< metal2 >>
rect -7990 1060 -220 1070
rect -7990 960 -350 1060
rect -250 960 -220 1060
rect -7990 950 -220 960
rect -7990 -6140 -7870 950
rect -6360 780 5220 800
rect -6360 700 5120 780
rect 5200 700 5220 780
rect -6360 680 5220 700
rect -6360 -740 -6240 680
rect -760 -220 7340 -200
rect -760 -300 2560 -220
rect 2620 -300 7340 -220
rect -760 -320 7340 -300
rect -760 -560 -640 -320
rect -760 -620 -740 -560
rect -660 -620 -640 -560
rect -760 -640 -640 -620
rect -360 -560 7340 -540
rect -360 -620 -340 -560
rect -260 -620 7340 -560
rect -360 -640 7340 -620
rect -6360 -820 -6340 -740
rect -6260 -820 -6240 -740
rect -6360 -840 -6240 -820
rect -800 -1020 -700 -1000
rect -800 -1080 -780 -1020
rect -720 -1080 -700 -1020
rect -800 -1380 -700 -1080
rect 80 -1020 180 -1000
rect 80 -1080 100 -1020
rect 160 -1080 180 -1020
rect 80 -1380 180 -1080
rect -800 -1440 -780 -1380
rect -720 -1440 100 -1380
rect 160 -1440 180 -1380
rect -800 -1460 180 -1440
rect -2160 -1580 -2060 -1540
rect 1460 -1580 1560 -1540
rect -2160 -1640 -2140 -1580
rect -2080 -1640 -2060 -1580
rect -2160 -1660 -2060 -1640
rect -3260 -2220 -2740 -2200
rect -3260 -2280 -3240 -2220
rect -3180 -2280 -2820 -2220
rect -2760 -2280 -2740 -2220
rect -3260 -2300 -2740 -2280
rect -2160 -2660 -2120 -1660
rect -2160 -2780 -2060 -2660
rect -940 -1600 -820 -1580
rect -940 -1660 -920 -1600
rect -840 -1660 -820 -1600
rect -940 -1960 -820 -1660
rect -940 -2020 -920 -1960
rect -840 -2020 -820 -1960
rect -940 -2300 -820 -2020
rect -940 -2360 -920 -2300
rect -840 -2360 -820 -2300
rect -940 -2660 -820 -2360
rect -940 -2720 -920 -2660
rect -840 -2720 -820 -2660
rect -940 -2740 -820 -2720
rect 220 -1600 340 -1580
rect 220 -1660 240 -1600
rect 320 -1660 340 -1600
rect 220 -1960 340 -1660
rect 220 -2020 240 -1960
rect 320 -2020 340 -1960
rect 220 -2300 340 -2020
rect 220 -2360 240 -2300
rect 320 -2360 340 -2300
rect 220 -2660 340 -2360
rect 220 -2720 240 -2660
rect 320 -2720 340 -2660
rect 220 -2740 340 -2720
rect 1460 -1640 1480 -1580
rect 1540 -1640 1560 -1580
rect 4080 -1560 4860 -1540
rect 4080 -1620 4100 -1560
rect 4160 -1620 4780 -1560
rect 4840 -1620 4860 -1560
rect 4080 -1640 4860 -1620
rect 1460 -1660 1560 -1640
rect 1520 -2660 1560 -1660
rect -700 -2780 -600 -2760
rect -700 -2840 -680 -2780
rect -620 -2800 -600 -2780
rect -100 -2780 0 -2760
rect 1460 -2780 1560 -2660
rect 5500 -2140 7340 -2040
rect -100 -2800 -80 -2780
rect -620 -2840 -80 -2800
rect -20 -2840 0 -2780
rect -700 -2860 0 -2840
rect 5500 -2840 5600 -2140
rect 6150 -2220 6940 -2200
rect 6150 -2280 6170 -2220
rect 6230 -2280 6940 -2220
rect 6150 -2300 6940 -2280
rect 5500 -2900 5520 -2840
rect 5580 -2900 5600 -2840
rect 5500 -2920 5600 -2900
rect -1880 -2940 5600 -2920
rect -1880 -3000 -1860 -2940
rect -1800 -3000 5600 -2940
rect -1880 -3020 5600 -3000
rect 6470 -2840 6570 -2820
rect 6470 -2900 6490 -2840
rect 6550 -2900 6570 -2840
rect -5080 -3120 6020 -3100
rect -5080 -3180 -5060 -3120
rect -5000 -3180 2340 -3120
rect 2400 -3180 6020 -3120
rect -5080 -3200 6020 -3180
rect 5920 -3420 6020 -3200
rect 6470 -3420 6570 -2900
rect 5920 -3520 6570 -3420
rect 6780 -3680 6940 -2300
rect 6500 -3840 6940 -3680
rect 4420 -3960 6220 -3940
rect 4420 -4020 4460 -3960
rect 4520 -4020 6120 -3960
rect 6180 -4020 6220 -3960
rect 4420 -4040 6220 -4020
rect -7990 -6160 -7020 -6140
rect -7990 -6280 -7160 -6160
rect -7040 -6280 -7020 -6160
rect -7990 -6300 -7020 -6280
rect 6500 -62720 6660 -3840
rect 6500 -62800 6540 -62720
rect 6620 -62800 6660 -62720
rect 6500 -62840 6660 -62800
<< via2 >>
rect -2120 -2660 -2060 -1660
rect -920 -1660 -840 -1600
rect -920 -2020 -840 -1960
rect -920 -2360 -840 -2300
rect -920 -2720 -840 -2660
rect 240 -1660 320 -1600
rect 240 -2020 320 -1960
rect 240 -2360 320 -2300
rect 240 -2720 320 -2660
rect 1460 -2660 1520 -1660
<< mimcap >>
rect -2130 -1740 -1130 -1660
rect -2130 -2580 -2050 -1740
rect -1210 -2580 -1130 -1740
rect -2130 -2660 -1130 -2580
rect 530 -1740 1530 -1660
rect 530 -2580 610 -1740
rect 1450 -2580 1530 -1740
rect 530 -2660 1530 -2580
<< mimcapcontact >>
rect -2050 -2580 -1210 -1740
rect 610 -2580 1450 -1740
<< metal3 >>
rect -2160 -1660 -2060 -1540
rect -2160 -2660 -2120 -1660
rect -2160 -2780 -2060 -2660
rect -940 -1600 -820 -1580
rect -940 -1660 -920 -1600
rect -840 -1660 -820 -1600
rect -940 -1960 -820 -1660
rect -940 -2020 -920 -1960
rect -840 -2020 -820 -1960
rect -940 -2300 -820 -2020
rect -940 -2360 -920 -2300
rect -840 -2360 -820 -2300
rect -940 -2660 -820 -2360
rect -940 -2720 -920 -2660
rect -840 -2720 -820 -2660
rect -940 -2740 -820 -2720
rect 220 -1600 340 -1580
rect 220 -1660 240 -1600
rect 320 -1660 340 -1600
rect 220 -1960 340 -1660
rect 220 -2020 240 -1960
rect 320 -2020 340 -1960
rect 220 -2300 340 -2020
rect 220 -2360 240 -2300
rect 320 -2360 340 -2300
rect 220 -2660 340 -2360
rect 220 -2720 240 -2660
rect 320 -2720 340 -2660
rect 220 -2740 340 -2720
rect 1460 -1660 1560 -1540
rect 1520 -2660 1560 -1660
rect 1460 -2780 1560 -2660
<< via3 >>
rect -920 -1660 -840 -1600
rect -920 -2020 -840 -1960
rect -920 -2360 -840 -2300
rect -920 -2720 -840 -2660
rect 240 -1660 320 -1600
rect 240 -2020 320 -1960
rect 240 -2360 320 -2300
rect 240 -2720 320 -2660
<< metal4 >>
rect -2250 -1600 -770 -1540
rect -2250 -1660 -920 -1600
rect -840 -1607 -770 -1600
rect -2250 -2660 -2130 -1660
rect -1130 -2660 -920 -1660
rect -2250 -2720 -920 -2660
rect -832 -2713 -770 -1607
rect -840 -2720 -770 -2713
rect -2250 -2780 -770 -2720
rect 170 -1600 1650 -1540
rect 170 -1607 240 -1600
rect 170 -2713 232 -1607
rect 320 -1660 1650 -1600
rect 320 -2660 530 -1660
rect 1530 -2660 1650 -1660
rect 170 -2720 240 -2713
rect 320 -2720 1650 -2660
rect 170 -2780 1650 -2720
<< via4 >>
rect -920 -1660 -840 -1607
rect -840 -1660 -832 -1607
rect -920 -1960 -832 -1660
rect -920 -2020 -840 -1960
rect -840 -2020 -832 -1960
rect -920 -2300 -832 -2020
rect -920 -2360 -840 -2300
rect -840 -2360 -832 -2300
rect -920 -2660 -832 -2360
rect -920 -2713 -840 -2660
rect -840 -2713 -832 -2660
rect 232 -1660 240 -1607
rect 240 -1660 320 -1607
rect 232 -1960 320 -1660
rect 232 -2020 240 -1960
rect 240 -2020 320 -1960
rect 232 -2300 320 -2020
rect 232 -2360 240 -2300
rect 240 -2360 320 -2300
rect 232 -2660 320 -2360
rect 232 -2713 240 -2660
rect 240 -2713 320 -2660
<< metal5 >>
rect -920 -1607 -832 -1597
rect -920 -2723 -832 -2713
rect 232 -1607 320 -1597
rect 232 -2723 320 -2713
use cap_mim_2p0fF_ZHL43H  cap_mim_2p0fF_ZHL43H_0
timestamp 1757657021
transform 1 0 -1510 0 1 -2160
box -740 -620 740 620
use cap_mim_2p0fF_ZHL43H  cap_mim_2p0fF_ZHL43H_2
timestamp 1757657021
transform -1 0 910 0 1 -2160
box -740 -620 740 620
use nfet_03v3_EF5H4U  nfet_03v3_EF5H4U_1
timestamp 1757524825
transform 1 0 6290 0 1 -3184
box -140 -156 140 156
use nfet_03v3_N5W335  nfet_03v3_N5W335_2
timestamp 1757529591
transform 1 0 -1440 0 1 -32928
box -140 -852 140 852
use nfet_03v3_N5WHL5  nfet_03v3_N5WHL5_1
timestamp 1757529591
transform 1 0 5560 0 1 -32228
box -140 -152 140 152
use nfet_03v3_NL3C35  nfet_03v3_NL3C35_1
timestamp 1757529591
transform 1 0 -4640 0 1 -32540
box -140 -460 140 460
use nfet_03v3_NL3C35  nfet_03v3_NL3C35_2
timestamp 1757529591
transform 1 0 -6240 0 1 -32540
box -140 -460 140 460
use nfet_03v3_NL3C35  nfet_03v3_NL3C35_3
timestamp 1757529591
transform 1 0 -5440 0 1 -32540
box -140 -460 140 460
use nfet_03v3_NMLPX4  nfet_03v3_NMLPX4_1
timestamp 1757063525
transform 0 1 -3132 -1 0 -1220
box -140 -2308 140 2308
use nfet_03v3_NMLPX4  nfet_03v3_NMLPX4_2
timestamp 1757063525
transform 0 1 2548 -1 0 -1220
box -140 -2308 140 2308
use nfet_03v3_NP3335  nfet_03v3_NP3335_0
timestamp 1757535309
transform 0 1 -5032 -1 0 -2060
box -140 -1748 140 1748
use nfet_03v3_NP3335  nfet_03v3_NP3335_1
timestamp 1757535309
transform 0 1 -5032 -1 0 -2440
box -140 -1748 140 1748
use nfet_03v3_NPKKZ4  nfet_03v3_NPKKZ4_1
timestamp 1757527981
transform 1 0 1560 0 1 -32432
box -140 -348 140 348
use nfet_03v3_NPKKZ4  nfet_03v3_NPKKZ4_2
timestamp 1757527981
transform 1 0 2360 0 1 -32432
box -140 -348 140 348
use nfet_03v3_NPKKZ4  nfet_03v3_NPKKZ4_3
timestamp 1757527981
transform 1 0 3160 0 1 -32432
box -140 -348 140 348
use nfet_03v3_NPKKZ4  nfet_03v3_NPKKZ4_4
timestamp 1757527981
transform 1 0 3960 0 1 -32432
box -140 -348 140 348
use nfet_03v3_NPKKZ4  nfet_03v3_NPKKZ4_5
timestamp 1757527981
transform 1 0 760 0 1 -32432
box -140 -348 140 348
use nfet_03v3_NUG935  nfet_03v3_NUG935_0
timestamp 1757012598
transform 0 1 -4252 -1 0 -780
box -140 -1188 140 1188
use nfet_03v3_NUG935  nfet_03v3_NUG935_1
timestamp 1757012598
transform 0 1 -1792 -1 0 -780
box -140 -1188 140 1188
use nfet_03v3_NUG935  nfet_03v3_NUG935_2
timestamp 1757012598
transform 0 1 3668 -1 0 -780
box -140 -1188 140 1188
use nfet_03v3_NUG935  nfet_03v3_NUG935_3
timestamp 1757012598
transform 0 1 1168 -1 0 -780
box -140 -1188 140 1188
use pfet_03v3_6ZJ338  pfet_03v3_6ZJ338_1
timestamp 1757524825
transform 1 0 6292 0 1 -2522
box -202 -218 202 218
use pplus_u_CRD77H  pplus_u_CRD77H_0
timestamp 1757010180
transform 0 -1 712 1 0 166
box -286 -772 286 772
use pplus_u_CRD77H  pplus_u_CRD77H_2
timestamp 1757010180
transform 0 -1 -1308 1 0 166
box -286 -772 286 772
use ppolyf_s_LGHZ3Z  ppolyf_s_LGHZ3Z_0
timestamp 1757698756
transform 0 1 6169 -1 0 -1222
box -258 -789 258 789
use ppolyf_s_LGHZ3Z  ppolyf_s_LGHZ3Z_1
timestamp 1757698756
transform 0 1 -6951 -1 0 -1222
box -258 -789 258 789
use ppolyf_u_1k_4GNJYW  ppolyf_u_1k_4GNJYW_1
timestamp 1757535624
transform 1 0 -7104 0 1 -4332
box -336 -1108 336 1108
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_0
timestamp 1757065516
transform 1 0 756 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_1
timestamp 1757065516
transform 1 0 1556 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_2
timestamp 1757065516
transform 1 0 2356 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_3
timestamp 1757065516
transform 1 0 3156 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_4
timestamp 1757065516
transform 1 0 3956 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_5
timestamp 1757065516
transform 1 0 5556 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_6
timestamp 1757065516
transform 1 0 -1444 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_7
timestamp 1757065516
transform 1 0 -2244 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_8
timestamp 1757065516
transform 1 0 -3844 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_9
timestamp 1757065516
transform 1 0 -5444 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_10
timestamp 1757065516
transform 1 0 -6244 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_11
timestamp 1757065516
transform 1 0 -4644 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_12
timestamp 1757065516
transform 1 0 -2244 0 1 -48282
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_13
timestamp 1757065516
transform 1 0 -1444 0 1 -48282
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_14
timestamp 1757065516
transform 1 0 756 0 1 -48242
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_15
timestamp 1757065516
transform 1 0 1556 0 1 -48242
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_16
timestamp 1757065516
transform 1 0 2356 0 1 -48242
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_17
timestamp 1757065516
transform 1 0 3156 0 1 -48242
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_18
timestamp 1757065516
transform 1 0 3956 0 1 -48242
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_19
timestamp 1757065516
transform 1 0 5556 0 1 -48242
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_20
timestamp 1757065516
transform 1 0 -3844 0 1 -48282
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_21
timestamp 1757065516
transform 1 0 -4644 0 1 -48282
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_22
timestamp 1757065516
transform 1 0 -5444 0 1 -48282
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_23
timestamp 1757065516
transform 1 0 -6244 0 1 -48282
box -336 -14358 336 14358
<< labels >>
rlabel metal1 7320 -4040 7420 -3940 1 AGND
rlabel metal1 7220 -1280 7340 -1160 1 RF-
rlabel metal1 -8260 -500 -8140 -380 1 IF+
rlabel metal1 -380 1360 -220 1520 1 VDD
rlabel metal1 7220 -840 7340 -720 1 LO+
rlabel metal2 7240 -640 7340 -540 1 LO-
rlabel metal2 7220 -320 7340 -200 1 IF-
rlabel metal1 -8260 -1280 -8140 -1160 1 RF+
rlabel metal1 7180 -1940 7340 -1780 1 MOSBIUS
rlabel metal2 7240 -2140 7340 -2040 1 VINSwitch
<< end >>
